--
--  File Name:         PcieContext.vhd
--  Design Unit Name:  PcieContext
--  Revision:          OSVVM MODELS STANDARD VERSION
--
--  Maintainer:        Simon Southwell      email:  simon.southwell@gmail.com
--  Contributor(s):
--     Simon Southwell      simon.southwell@gmail.com
--
--
--  Description:
--      Pcie GEN1/2 model
--
--  Revision History:
--    Date      Version    Description
--    07/2025   2026.01    Initial version
--
--
--  This file is part of OSVVM.
--
--  Copyright (c) 2025 by [OSVVM Authors](../../AUTHORS.md).
--
--  Licensed under the Apache License, Version 2.0 (the "License") ;
--  you may not use this file except in compliance with the License.
--  You may obtain a copy of the License at
--
--      https://www.apache.org/licenses/LICENSE-2.0
--
--  Unless required by applicable law or agreed to in writing, software
--  distributed under the License is distributed on an "AS IS" BASIS,
--  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--  See the License for the specific language governing permissions and
--  limitations under the License.
--
context PcieContext is

    library osvvm_common ;
    context osvvm_common.OsvvmCommonContext ;

    library osvvm_pcie ;

    use osvvm_pcie.PcieInterfacePkg.all ;
    use osvvm_pcie.PcieOptionsPkg.all ;
    use osvvm_pcie.PcieComponentPkg.all ;

end context PcieContext ;